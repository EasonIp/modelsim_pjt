`timescale 1ns/1ns
`define tp 1
module block_nonblock(Clk,Rst_n,a,b,c,out);

	input Clk;
	input Rst_n;
	input a,b,c;
	output reg [1:0]out;
	
	//out = a + b + c;
	
	//d = a+b;
	//out = d + c;
	
	reg [1:0] d;
	
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		out <= 2'b0;
	else begin
		out <= a + b + c;
	end
	
endmodule
