library ieee;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use ieee.std_logic_1164.all;
ENTITY sinb IS 
    PORT( CLK:IN STD_LOGIC;
          dout:OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END;

ARCHITECTURE arch OF sinb IS
  signal q1: integer range 0 to 400;
  signal dat: integer range -200 to 200;
  BEGIN
   PROCESS(CLK)
      BEGIN
       IF CLK'EVENT AND CLK='1' THEN 
          if q1=399 then  
               q1<=0;
          else 
               q1<=q1+1;
          end if;
case q1 is
when    0=>dat<=-200;
when    1=>dat<=-200;
when    2=>dat<=-200;
when    3=>dat<=-200;
when    4=>dat<=-200;
when    5=>dat<=-200;
when    6=>dat<=-200;
when    7=>dat<=-199;
when    8=>dat<=-199;
when    9=>dat<=-199;
when    10=>dat<=-198;
when    11=>dat<=-198;
when    12=>dat<=-197;
when    13=>dat<=-196;
when    14=>dat<=-196;
when    15=>dat<=-195;
when    16=>dat<=-194;
when    17=>dat<=-193;
when    18=>dat<=-193;
when    19=>dat<=-192;
when    20=>dat<=-191;
when    21=>dat<=-190;
when    22=>dat<=-189;
when    23=>dat<=-188;
when    24=>dat<=-186;
when    25=>dat<=-185;
when    26=>dat<=-184;
when    27=>dat<=-183;
when    28=>dat<=-181;
when    29=>dat<=-180;
when    30=>dat<=-179;
when    31=>dat<=-177;
when    32=>dat<=-176;
when    33=>dat<=-174;
when    34=>dat<=-173;
when    35=>dat<=-171;
when    36=>dat<=-169;
when    37=>dat<=-168;
when    38=>dat<=-166;
when    39=>dat<=-164;
when    40=>dat<=-162;
when    41=>dat<=-160;
when    42=>dat<=-159;
when    43=>dat<=-157;
when    44=>dat<=-155;
when    45=>dat<=-153;
when    46=>dat<=-151;
when    47=>dat<=-148;
when    48=>dat<=-146;
when    49=>dat<=-144;
when    50=>dat<=-142;
when    51=>dat<=-140;
when    52=>dat<=-137;
when    53=>dat<=-135;
when    54=>dat<=-133;
when    55=>dat<=-130;
when    56=>dat<=-128;
when    57=>dat<=-126;
when    58=>dat<=-123;
when    59=>dat<=-121;
when    60=>dat<=-118;
when    61=>dat<=-116;
when    62=>dat<=-113;
when    63=>dat<=-110;
when    64=>dat<=-108;
when    65=>dat<=-105;
when    66=>dat<=-102;
when    67=>dat<=-100;
when    68=>dat<=-97;
when    69=>dat<=-94;
when    70=>dat<=-91;
when    71=>dat<=-88;
when    72=>dat<=-86;
when    73=>dat<=-83;
when    74=>dat<=-80;
when    75=>dat<=-77;
when    76=>dat<=-74;
when    77=>dat<=-71;
when    78=>dat<=-68;
when    79=>dat<=-65;
when    80=>dat<=-62;
when    81=>dat<=-59;
when    82=>dat<=-56;
when    83=>dat<=-53;
when    84=>dat<=-50;
when    85=>dat<=-47;
when    86=>dat<=-44;
when    87=>dat<=-41;
when    88=>dat<=-38;
when    89=>dat<=-35;
when    90=>dat<=-32;
when    91=>dat<=-29;
when    92=>dat<=-26;
when    93=>dat<=-22;
when    94=>dat<=-19;
when    95=>dat<=-16;
when    96=>dat<=-13;
when    97=>dat<=-10;
when    98=>dat<=-7;
when    99=>dat<=-4;
when    100=>dat<=0;
when    101=>dat<=3;
when    102=>dat<=6;
when    103=>dat<=9;
when    104=>dat<=12;
when    105=>dat<=15;
when    106=>dat<=18;
when    107=>dat<=21;
when    108=>dat<=25;
when    109=>dat<=28;
when    110=>dat<=31;
when    111=>dat<=34;
when    112=>dat<=37;
when    113=>dat<=40;
when    114=>dat<=43;
when    115=>dat<=46;
when    116=>dat<=49;
when    117=>dat<=52;
when    118=>dat<=55;
when    119=>dat<=58;
when    120=>dat<=61;
when    121=>dat<=64;
when    122=>dat<=67;
when    123=>dat<=70;
when    124=>dat<=73;
when    125=>dat<=76;
when    126=>dat<=79;
when    127=>dat<=82;
when    128=>dat<=85;
when    129=>dat<=87;
when    130=>dat<=90;
when    131=>dat<=93;
when    132=>dat<=96;
when    133=>dat<=99;
when    134=>dat<=101;
when    135=>dat<=104;
when    136=>dat<=107;
when    137=>dat<=109;
when    138=>dat<=112;
when    139=>dat<=115;
when    140=>dat<=117;
when    141=>dat<=120;
when    142=>dat<=122;
when    143=>dat<=125;
when    144=>dat<=127;
when    145=>dat<=129;
when    146=>dat<=132;
when    147=>dat<=134;
when    148=>dat<=136;
when    149=>dat<=139;
when    150=>dat<=141;
when    151=>dat<=143;
when    152=>dat<=145;
when    153=>dat<=147;
when    154=>dat<=150;
when    155=>dat<=152;
when    156=>dat<=154;
when    157=>dat<=156;
when    158=>dat<=158;
when    159=>dat<=159;
when    160=>dat<=161;
when    161=>dat<=163;
when    162=>dat<=165;
when    163=>dat<=167;
when    164=>dat<=168;
when    165=>dat<=170;
when    166=>dat<=172;
when    167=>dat<=173;
when    168=>dat<=175;
when    169=>dat<=176;
when    170=>dat<=178;
when    171=>dat<=179;
when    172=>dat<=180;
when    173=>dat<=182;
when    174=>dat<=183;
when    175=>dat<=184;
when    176=>dat<=185;
when    177=>dat<=187;
when    178=>dat<=188;
when    179=>dat<=189;
when    180=>dat<=190;
when    181=>dat<=191;
when    182=>dat<=192;
when    183=>dat<=192;
when    184=>dat<=193;
when    185=>dat<=194;
when    186=>dat<=195;
when    187=>dat<=195;
when    188=>dat<=196;
when    189=>dat<=197;
when    190=>dat<=197;
when    191=>dat<=198;
when    192=>dat<=198;
when    193=>dat<=198;
when    194=>dat<=199;
when    195=>dat<=199;
when    196=>dat<=199;
when    197=>dat<=199;
when    198=>dat<=199;
when    199=>dat<=199;
when    200=>dat<=200;
when    201=>dat<=199;
when    202=>dat<=199;
when    203=>dat<=199;
when    204=>dat<=199;
when    205=>dat<=199;
when    206=>dat<=199;
when    207=>dat<=198;
when    208=>dat<=198;
when    209=>dat<=198;
when    210=>dat<=197;
when    211=>dat<=197;
when    212=>dat<=196;
when    213=>dat<=195;
when    214=>dat<=195;
when    215=>dat<=194;
when    216=>dat<=193;
when    217=>dat<=192;
when    218=>dat<=192;
when    219=>dat<=191;
when    220=>dat<=190;
when    221=>dat<=189;
when    222=>dat<=188;
when    223=>dat<=187;
when    224=>dat<=185;
when    225=>dat<=184;
when    226=>dat<=183;
when    227=>dat<=182;
when    228=>dat<=180;
when    229=>dat<=179;
when    230=>dat<=178;
when    231=>dat<=176;
when    232=>dat<=175;
when    233=>dat<=173;
when    234=>dat<=172;
when    235=>dat<=170;
when    236=>dat<=168;
when    237=>dat<=167;
when    238=>dat<=165;
when    239=>dat<=163;
when    240=>dat<=161;
when    241=>dat<=159;
when    242=>dat<=158;
when    243=>dat<=156;
when    244=>dat<=154;
when    245=>dat<=152;
when    246=>dat<=150;
when    247=>dat<=147;
when    248=>dat<=145;
when    249=>dat<=143;
when    250=>dat<=141;
when    251=>dat<=139;
when    252=>dat<=136;
when    253=>dat<=134;
when    254=>dat<=132;
when    255=>dat<=129;
when    256=>dat<=127;
when    257=>dat<=125;
when    258=>dat<=122;
when    259=>dat<=120;
when    260=>dat<=117;
when    261=>dat<=115;
when    262=>dat<=112;
when    263=>dat<=109;
when    264=>dat<=107;
when    265=>dat<=104;
when    266=>dat<=101;
when    267=>dat<=99;
when    268=>dat<=96;
when    269=>dat<=93;
when    270=>dat<=90;
when    271=>dat<=87;
when    272=>dat<=85;
when    273=>dat<=82;
when    274=>dat<=79;
when    275=>dat<=76;
when    276=>dat<=73;
when    277=>dat<=70;
when    278=>dat<=67;
when    279=>dat<=64;
when    280=>dat<=61;
when    281=>dat<=58;
when    282=>dat<=55;
when    283=>dat<=52;
when    284=>dat<=49;
when    285=>dat<=46;
when    286=>dat<=43;
when    287=>dat<=40;
when    288=>dat<=37;
when    289=>dat<=34;
when    290=>dat<=31;
when    291=>dat<=28;
when    292=>dat<=25;
when    293=>dat<=21;
when    294=>dat<=18;
when    295=>dat<=15;
when    296=>dat<=12;
when    297=>dat<=9;
when    298=>dat<=6;
when    299=>dat<=3;
when    300=>dat<=0;
when    301=>dat<=-4;
when    302=>dat<=-7;
when    303=>dat<=-10;
when    304=>dat<=-13;
when    305=>dat<=-16;
when    306=>dat<=-19;
when    307=>dat<=-22;
when    308=>dat<=-26;
when    309=>dat<=-29;
when    310=>dat<=-32;
when    311=>dat<=-35;
when    312=>dat<=-38;
when    313=>dat<=-41;
when    314=>dat<=-44;
when    315=>dat<=-47;
when    316=>dat<=-50;
when    317=>dat<=-53;
when    318=>dat<=-56;
when    319=>dat<=-59;
when    320=>dat<=-62;
when    321=>dat<=-65;
when    322=>dat<=-68;
when    323=>dat<=-71;
when    324=>dat<=-74;
when    325=>dat<=-77;
when    326=>dat<=-80;
when    327=>dat<=-83;
when    328=>dat<=-86;
when    329=>dat<=-88;
when    330=>dat<=-91;
when    331=>dat<=-94;
when    332=>dat<=-97;
when    333=>dat<=-100;
when    334=>dat<=-102;
when    335=>dat<=-105;
when    336=>dat<=-108;
when    337=>dat<=-110;
when    338=>dat<=-113;
when    339=>dat<=-116;
when    340=>dat<=-118;
when    341=>dat<=-121;
when    342=>dat<=-123;
when    343=>dat<=-126;
when    344=>dat<=-128;
when    345=>dat<=-130;
when    346=>dat<=-133;
when    347=>dat<=-135;
when    348=>dat<=-137;
when    349=>dat<=-140;
when    350=>dat<=-142;
when    351=>dat<=-144;
when    352=>dat<=-146;
when    353=>dat<=-148;
when    354=>dat<=-151;
when    355=>dat<=-153;
when    356=>dat<=-155;
when    357=>dat<=-157;
when    358=>dat<=-159;
when    359=>dat<=-160;
when    360=>dat<=-162;
when    361=>dat<=-164;
when    362=>dat<=-166;
when    363=>dat<=-168;
when    364=>dat<=-169;
when    365=>dat<=-171;
when    366=>dat<=-173;
when    367=>dat<=-174;
when    368=>dat<=-176;
when    369=>dat<=-177;
when    370=>dat<=-179;
when    371=>dat<=-180;
when    372=>dat<=-181;
when    373=>dat<=-183;
when    374=>dat<=-184;
when    375=>dat<=-185;
when    376=>dat<=-186;
when    377=>dat<=-188;
when    378=>dat<=-189;
when    379=>dat<=-190;
when    380=>dat<=-191;
when    381=>dat<=-192;
when    382=>dat<=-193;
when    383=>dat<=-193;
when    384=>dat<=-194;
when    385=>dat<=-195;
when    386=>dat<=-196;
when    387=>dat<=-196;
when    388=>dat<=-197;
when    389=>dat<=-198;
when    390=>dat<=-198;
when    391=>dat<=-199;
when    392=>dat<=-199;
when    393=>dat<=-199;
when    394=>dat<=-200;
when    395=>dat<=-200;
when    396=>dat<=-200;
when    397=>dat<=-200;
when    398=>dat<=-200;
when    399=>dat<=-200;



when   others=> dat<=0;
end case;
 dout<= conv_std_logic_vector (dat,16);
END IF;
 
  
   END PROCESS;
END;
